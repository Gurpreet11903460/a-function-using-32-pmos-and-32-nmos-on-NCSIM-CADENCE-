module functionpmos(a,b,c,d,y);
input a,b,c,d;
output y;
supply1 vdd;
supply0 vss;
wire abar,bbar,cbar,dbar,w1,w2,w3,w4,w5,w6,w7,w8;
wire w9,w10,w11,w12,w13,w14,w15,w16,w17,w18,w19,w20,w21,w22,w23;
wire w24,w25,w26,w27,w28,w29,w30,w31,w32;
not n89(abar,a);
not n77(bbar,b);
not n33(cbar,c);
not n44(dbar,d);
pmos p1(w1,vdd,abar);
pmos p2(w1,vdd,bbar);
pmos p3(w1,vdd,cbar);
pmos p4(w1,vdd,dbar);
pmos p5(w2,w1,abar);
pmos p6(w2,w1,bbar);
pmos p7(w2,w1,c);
pmos p8(w2,w1,dbar);
pmos p9(w3,w2,abar);
pmos p10(w3,w2,bbar);
pmos p11(w3,w2,c);
pmos p12(w3,w2,d);
pmos p13(w4,w3,abar);
pmos p14(w4,w3,b);
pmos p15(w4,w3,c);
pmos p16(w4,w3,dbar);
pmos p17(w5,w4,abar);
pmos p18(w5,w4,b);
pmos p19(w5,w4,c);
pmos p20(w5,w4,d);
pmos p21(w6,w5,a);
pmos p22(w6,w5,bbar);
pmos p23(w6,w5,c);
pmos p24(w6,w5,dbar);
pmos p25(w7,w6,a);
pmos p26(w7,w6,b);
pmos p27(w7,w6,cbar);
pmos p28(w7,w6,dbar);
pmos p29(w8,w7,a);
pmos p30(w8,w7,b);
pmos p31(w8,w7,cbar);
pmos p32(w8,w7,d);
nmos n1(w8,w9,abar);
nmos n2(w9,w10,bbar);
nmos n3(w10,w11,cbar);
nmos n4(w11,vss,dbar);
nmos n5(w8,w12,abar);
nmos n6(w12,w13,bbar);
nmos n7(w13,w14,c);
nmos n8(w14,vss,dbar);
nmos n9(w8,w15,abar);
nmos n10(w15,w16,bbar);
nmos n11(w16,w17,c);
nmos n12(w17,vss,d);
nmos n13(w8,w18,abar);
nmos n14(w18,w19,b);
nmos n15(w19,w20,c);
nmos n16(w20,vss,dbar);
nmos n17(w8,w21,abar);
nmos n18(w21,w22,b);
nmos n19(w22,w23,c);
nmos n20(w23,vss,d);
nmos n21(w8,w24,a);
nmos n22(w24,w25,bbar);
nmos n23(w25,w26,c);
nmos n24(w26,vss,dbar);
nmos n25(w8,w27,a);
nmos n26(w27,w28,b);
nmos n27(w28,w29,cbar);
nmos n28(w29,vss,dbar);
nmos n29(w8,w30,a);
nmos n30(w30,w31,b);
nmos n31(w31,w32,cbar);
nmos n32(w32,vss,d);
not n88(y,w8);
endmodule

module functionpmostb();
reg a,b,c,d;
wire y;
functionpmos f1(a,b,c,d,y);
initial
begin
a=0;b=0;c=0;d=0;
#2 a=0;b=0;c=0;d=1;
#2 a=0;b=0;c=1;d=0;
#2 a=0;b=0;c=1;d=1;
#2 a=0;b=1;c=0;d=0;
#2 a=0;b=1;c=0;d=1;
#2 a=0;b=1;c=1;d=0;
#2 a=0;b=1;c=1;d=1;
#2 a=1;b=0;c=0;d=0;
#2 a=1;b=0;c=0;d=1;
#2 a=1;b=0;c=1;d=0;
#2 a=1;b=0;c=1;d=1;
#2 a=1;b=1;c=0;d=0;
#2 a=1;b=1;c=0;d=1;
#2 a=1;b=1;c=1;d=0;
#2 a=1;b=1;c=1;d=1;
#2 $stop;
end
endmodule
